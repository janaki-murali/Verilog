module not_gate(
  input x,
  output y);
  assign y=~x;
endmodule
